// SPDX-License-Identifier: MIT

/* This file contains the frequently used defaults. */

/* ------------------------------------------------------------------------- */


/*
 * Word size for the processor.
 * This also defines the register file width, bus width, etc.
 */
`define WORD_SIZE       32
`define L2_WORD_SIZE    5   /* log2(WORD_SIZE) = Number of bits. */


/* Number of registers (as in x0-x31) in the register file. */
`define REG_FILE_SIZE       32
`define L2_REG_FILE_SIZE    5


/* ------------------------------------------------------------------------- */


/* End of file. */
