`include "core.pkg"

module core
  (
    input clk,
    input rst
  );
  
  
  
  
  
endmodule
